`define NO_OF_PACKETS 20
static int ERROR=0;