`define UART_IDLE 1
`define UART_START 0
`define UART_STOP 1

`define WORD_LENGTH 8
`define PARITY_LENGTH 1

`define COUNTER_START 1
`define COUNTER_STOP 0

`define Tx_BUSY 0
`define Tx_READY 1

`define Tx_CLKRATE 1_000_000
`define Rx_CLKRATE 1_000_000
`define BAUD 9600

`define PCKT_OK 0
`define PCKT_NOT_OK 1